/Users/karstenbecker/Dropbox/PSHDL/PSHDLCode/lib/pshdl_pkg.vhd